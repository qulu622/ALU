module MULTIPLIER( inputA, inputB, result, reset, clk, Signal);input reset,clk;input [31:0]inputA, inputB;input [5:0]Signal ;output [63:0]result;reg [63:0] MCAND ;reg [31:0] MLER ;reg [63:0] product;reg [5:0]count ;parameter MULTU = 6'd25;always @( Signal or inputA or inputB ) begin	if ( Signal == MULTU ) 	begin		count = 6'd0;		MCAND[63:0] = {32'b0,inputA} ;		MLER = inputB ;					product = 0 ;	endendalways @( posedge clk )begin	if(reset) 	begin 					product = 64'd0;	end	else if( count < 32 )	begin 		if( MLER[0] == 1'b1 )		begin 			product = product + MCAND ;		end		else 		begin			product = product;		end				MCAND = MCAND << 1 ;		MLER = MLER >> 1 ;		count = count + 6'd1 ;				endendassign result = product;endmodule